module HA(a,b,sum,carry );
input a,b;
output reg sum, carry;
  assign sum =a+b;
  assign carry=ab;
endmodule 
